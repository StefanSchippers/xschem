* comp3_read.cir

.subckt comp3_read PLUS OUT MINUS
v1 x 0 1.1
e1 out x plus minus 0.5
.ends
